package adapter_package;

        `include "adapter_env.sv"

endpackage